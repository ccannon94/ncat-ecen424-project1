library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity code_timeout_timer is
  port(enable, reset, clk : in std_logic; done : out std_logic);
end entity code_timeout_timer;

architecture code_timeout_behavior is

end architecture code_timeout_behavior;
